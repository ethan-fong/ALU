module part3(A,B,Function,ALUout);
	input [3:0]A;
	input [3:0]B;
	input [2:0]Function;
	output [7:0]ALUout;
	wire w0;
	wire [3:0]w1;
	wire [4:0]tmp;
	assign tmp = A+B;
	part2 forALU (A[3:0],B[3:0],1'b0,w1[3:0],w0);
	reg [7:0]ALUout;
		always @(*)
			begin
				case(Function[2:0])
					3'b000: ALUout[7:0]={3'b000,w0,w1[3:0]};
					3'b001: ALUout[7:0]={3'b000,tmp[4],tmp[3:0]}; //work in progress
					3'b010: ALUout[7:0]={B[3],B[3],B[3],B[3],B[3:0]};
					3'b011: ALUout[7:0]={7'b0000000,|{A[3:0],B[3:0]}};
					3'b100: ALUout[7:0]={7'b0000000,&{A[3:0],B[3:0]}};
					3'b101: ALUout[7:0]={A[3:0],B[3:0]};
					default: ALUout[7:0]=8'b11011110;
				endcase
			end
			
endmodule

module fulladder(bit_1,bit_2,c_in,c_out,s);
	input bit_1,bit_2,c_in;
	output c_out,s;
	assign s = bit_1^bit_2^c_in;
	assign c_out = (bit_1&bit_2)|(bit_1&c_in)|(bit_2&c_in);
endmodule

module hex_decoder (c,display);
	input  [3:0]c;
	output [6:0]display;
	assign display[0] = ~(((~c[0])&(~c[1])&(~c[2])&(~c[3])) 
|((~c[0])&(c[1])&(~c[2])&(~c[3])) |((~c[3])&(~c[2])&(c[1])&(c[0]))
|((~c[3])&(c[2])&(~c[1])&(c[0]))|((~c[3])&(c[2])&(c[1])&(~c[0]))
|((~c[3])&(c[2])&(c[1])&(c[0]))|((c[3])&(~c[2])&(~c[1])&(~c[0]))
|((c[3])&(~c[2])&(~c[1])&(c[0]))|((c[3])&(~c[2])&(c[1])&(~c[0]))
|((c[3])&(c[2])&(~c[1])&(~c[0]))|((c[3])&(c[2])&(c[1])&(~c[0]))|((c[3])&(c[2])&(c[1])&(c[0])));         

	assign display[1] =  ~(((~c[3])&(~c[2])&(~c[1])&(~c[0]))
 |((~c[3])&(~c[2])&(~c[1])&(c[0]))
 |((~c[3])&(~c[2])&(c[1])&(~c[0]))
 |((~c[3])&(~c[2])&(c[1])&(c[0])) 
|((~c[3])&(c[2])&(~c[1])&(~c[0]))
|((~c[3])&(c[2])&(c[1])&(c[0]))
|((c[3])&(~c[2])&(~c[1])&(~c[0]))
|((c[3])&(~c[2])&(~c[1])&(c[0]))
|((c[3])&(~c[2])&(c[1])&(~c[0]))
|((c[3])&(c[2])&(~c[1])&(c[0])));

assign display[2] =  ~(((~c[3])&(~c[2])&(~c[1])&(~c[0]))
 |((~c[3])&(~c[2])&(~c[1])&(c[0]))
 |((~c[3])&(~c[2])&(c[1])&(c[0])) 
|((~c[3])&(c[2])&(~c[1])&(~c[0]))
|((~c[3])&(c[2])&(~c[1])&(c[0]))
|((~c[3])&(c[2])&(c[1])&(~c[0]))
|((~c[3])&(c[2])&(c[1])&(c[0]))
|((c[3])&(~c[2])&(~c[1])&(~c[0]))
|((c[3])&(~c[2])&(~c[1])&(c[0]))
|((c[3])&(~c[2])&(c[1])&(~c[0]))
|((c[3])&(~c[2])&(c[1])&(c[0]))
|((c[3])&(c[2])&(~c[1])&(c[0])));

assign display[3] =  ~(((~c[3])&(~c[2])&(~c[1])&(~c[0]))
 |((~c[3])&(~c[2])&(c[1])&(~c[0]))
 |((~c[3])&(~c[2])&(c[1])&(c[0])) 
|((~c[3])&(c[2])&(~c[1])&(c[0]))
|((~c[3])&(c[2])&(c[1])&(~c[0]))
|((c[3])&(~c[2])&(~c[1])&(~c[0]))
|((c[3])&(~c[2])&(~c[1])&(c[0]))
|((c[3])&(~c[2])&(c[1])&(c[0]))
|((c[3])&(c[2])&(~c[1])&(~c[0]))
|((c[3])&(c[2])&(~c[1])&(c[0]))
|((c[3])&(c[2])&(c[1])&(~c[0])));

assign display[4] =  ~(((~c[3])&(~c[2])&(~c[1])&(~c[0]))
 |((~c[3])&(~c[2])&(c[1])&(~c[0]))
|((~c[3])&(c[2])&(c[1])&(~c[0]))
|((c[3])&(~c[2])&(~c[1])&(~c[0]))
|((c[3])&(~c[2])&(c[1])&(~c[0]))
|((c[3])&(~c[2])&(c[1])&(c[0]))
|((c[3])&(c[2])&(~c[1])&(~c[0]))
|((c[3])&(c[2])&(~c[1])&(c[0]))
|((c[3])&(c[2])&(c[1])&(~c[0]))
|((c[3])&(c[2])&(c[1])&(c[0])));        

assign display[5] =  ~(((~c[3])&(~c[2])&(~c[1])&(~c[0]))
|((~c[3])&(c[2])&(~c[1])&(~c[0]))
|((~c[3])&(c[2])&(~c[1])&(c[0]))
|((~c[3])&(c[2])&(c[1])&(~c[0]))
|((c[3])&(~c[2])&(~c[1])&(~c[0]))
|((c[3])&(~c[2])&(~c[1])&(c[0]))
|((c[3])&(~c[2])&(c[1])&(~c[0]))
|((c[3])&(~c[2])&(c[1])&(c[0]))
|((c[3])&(c[2])&(~c[1])&(~c[0]))
|((c[3])&(c[2])&(c[1])&(~c[0]))
|((c[3])&(c[2])&(c[1])&(c[0])));          

assign display[6] =  ~(((~c[3])&(~c[2])&(c[1])&(~c[0]))
 |((~c[3])&(~c[2])&(c[1])&(c[0])) 
|((~c[3])&(c[2])&(~c[1])&(~c[0]))
|((~c[3])&(c[2])&(~c[1])&(c[0]))
|((~c[3])&(c[2])&(c[1])&(~c[0]))
|((c[3])&(~c[2])&(~c[1])&(~c[0]))
|((c[3])&(~c[2])&(~c[1])&(c[0]))
|((c[3])&(~c[2])&(c[1])&(~c[0]))
|((c[3])&(~c[2])&(c[1])&(c[0]))
|((c[3])&(c[2])&(~c[1])&(c[0]))
|((c[3])&(c[2])&(c[1])&(~c[0]))
|((c[3])&(c[2])&(c[1])&(c[0])));

endmodule

module part2(a,b,c_in,s,c_out); //4 bit ripple adder
	input [3:0]a;
	input [3:0]b;
	input c_in;
	output [3:0]s;
	output c_out;
	wire w0,w1,w2,w3,w4;
	fulladder f1 (a[0],b[0],c_in,w0,s[0]);
	fulladder f2 (a[1],b[1],w0,w1,s[1]);
	fulladder f3 (a[2],b[2],w1,w2,s[2]);
	fulladder f4(a[3],b[3],w2,c_out,s[3]);
endmodule
